`timescale 1ns / 1ps
module Storage_filter_Mem(
    input re,we
    );

    reg [7:0] Mem [8:0];

endmodule

module dd (
    ports
);
    
endmodule
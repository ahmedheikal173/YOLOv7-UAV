`timescale 1ns / 1ps

module Padding_CBS_File(
    input clk,reset,count2_row_0,
    input [71:0] from_9_Reg,
    input [14:0]counter_Row,counter_Col,
    output reg [71:0] to_9_Reg
    );

    
        

endmodule

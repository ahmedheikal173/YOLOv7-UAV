module conv_FSM(img,filts,filtindex, mult_Loc_in,mult_Loc_out,free_mult_no, clk,rstn,en,     outdatimg,outdatflt);
//module conv_FSM(img,filts,filtindex, S,N,K, mult_Loc_in,mult_Loc_out,free_mult_no, clk,rstn,en,     outdatimg,outdatflt);
//moore fsm

//parameters
parameter IDLE = 3'b000;
parameter START = 3'b001;
parameter flt_ass = 3'b010;
parameter mult_ass = 3'b011;
parameter EXECUTE_full = 3'b100;
parameter EXECUTE_partial = 3'b101;
parameter READY = 3'b110;
parameter N = 32;
parameter F = 3;
parameter NF = 3;
parameter K=3;
parameter P=1;
parameter S=1;
parameter Nmult = 64; parameter Mmult = 6;
parameter W=64;


//input ports
//input [1:0] S,K; // ya2ema 1 aw 3
//input [63:0] N; // mesh aref a3melo kam lessa

input [Nmult-1:0] mult_Loc_in; // 0 free, 1 occupied
output reg [Nmult-1:0] mult_Loc_out; // 0 free, 1 occupied
input [Mmult-1:0] free_mult_no;
input [NF-1:0] filtindex;
input [W-1:0] filts [F-1:0][F-1:0][K-1:0];
input [W-1:0] img [N-1:0][N-1:0][K-1:0];
//input [W-1:0] filts [F*F*K-1:0];
//input [W-1:0] img [N*N*K-1:0];
input clk,rstn,en;


//output ports
output reg [W-1:0] outdatimg [N-1:0][N-1:0][K-1:0];
output reg [W-1:0] outdatflt [F-1:0][F-1:0][K-1:0];


// state regs
integer out_size,need_mults,i,j,k,iflt,jflt,kflt, ii,jj;
reg [2:0] cs,ns;

assign out_size = (N-F+2*P)/S +1;
assign need_mults = out_size*out_size*NF;
// next state logic
always@(*) begin
    case (cs)
        IDLE:
            begin
            
            
            end
        START:
            begin
                if (!en)
                    ns=IDLE;

            end
        flt_ass:
            begin
                if (!en)
                    ns=IDLE;

            end
        mult_ass://TODO:///////////////////////////////////////////////////////////////////
            begin
                // if (!en)
                //     ns=IDLE;
                // if (free_mult_no>=need_mults) begin
                //     // select free mults (FULL)
                //     for(k=0; k<K; k=k+1) begin
                //         for(j=0; j<N; j=j+S) begin
                //             for(i=0; i<N; i=i+S) begin
                //                 for (jflt=0,jflt<F,jflt=jflt+1)begin
                //                     for(iflt=0,iflt<F,iflt=iflt+1) begin
                //                         outdatimg = 
                //                     end
                //                 end
                //             end
                //         end
                //     end
                    
                // end
                // else begin
                //     //select free mults (PARTIAL)
                // end
            end
        EXECUTE_full:
            begin
                if (!en)
                    ns=IDLE;
                //for () begin


                //end

            end
        EXECUTE_partial:
            begin
                if (!en)
                    ns=IDLE;

            end
        READY:
            begin
                if (!en)
                    ns=IDLE;
                
            end
        default:
            begin
                ns=IDLE;
            end
    endcase    


end





///////////////////////////////

// state memory
always @ (posedge clk, negedge rstn) begin
    if (!rstn) begin
        cs <= IDLE;
    end
    else begin
        cs<=ns;
    end
end
////////////////////////////////


// output logic
always @(*) begin
    if (cs==IDLE) begin
    end
    if (cs==START) begin
    end
    if (cs==flt_ass) begin
    end
    if (cs==mult_ass) begin
        if (!en)
            ns=IDLE;
        if (free_mult_no>=need_mults) begin
            // select free mults (FULL)
            jj=0;
            for (ii=0;ii<Nmult;ii=ii+1) begin
                if (mult_Loc_in==0) begin
                    mult_Loc_out[jj]=mult_Loc_in[ii];
                    jj=jj+1;
                end
            end
            for(k=0; k<K; k=k+1) begin
                for(j=0; j<N; j=j+S) begin
                    for(i=0; i<N; i=i+S) begin
                        // for (ii=0;ii<Nmult;ii=ii+1) begin
                        //     if (mult_Loc_in==0) begin
                        //         mult_Loc_out[jj]=mult_Loc_in[ii];
                        //         jj=jj+1;
                        //     end
                        // end
                        for (kflt=0;kflt<F;kflt=kflt+1) begin
                            for(jflt=0;jflt<F;jflt=jflt+1) begin
                                for (iflt=0;iflt<F;iflt=iflt+1) begin
                                    outdatimg[i][j][k] = img [i][j][k];
                                    outdatflt[iflt][jflt][kflt] = filts[iflt][jflt][kflt];//TODO:///////////////////////////////////
                                    //outdatimg = img [i][j][k];
                                    //outdatflt = filts[iflt][jflt][kflt];//TODO:///////////////////////////////////
                                end
                            end
                        end
                    end
                end
            end
        end
        else begin
            //select free mults (PARTIAL)
            jj=0;
            for(k=0; k<K; k=k+1) begin
                for(j=0; j<N; j=j+S) begin
                    for(i=0; i<N; i=i+S) begin
                        for (ii=0;ii<Nmult;ii=ii+1) begin
                            if (mult_Loc_in==1) begin
                                mult_Loc_out[jj]=mult_Loc_in[ii];
                                jj=jj+1;
                            end
                        end
                        for (kflt=0;kflt<F;kflt=kflt+1) begin
                            for(jflt=0;jflt<F;jflt=jflt+1) begin
                                for (iflt=0;iflt<F;iflt=iflt+1) begin
                                    outdatimg[i][j][k] = img [i][j][k];
                                    outdatflt[iflt][jflt][kflt] = filts[iflt][jflt][kflt];//TODO:///////////////////////////////////
                                    //outdatimg = img [i][j][k];
                                    //outdatflt = filts[iflt][jflt][kflt];//TODO:///////////////////////////////////
                                end
                            end
                        end
                    end
                end
            end
        end
    end
    if (cs==EXECUTE_full) begin
    end
    if (cs==EXECUTE_partial) begin
    end
    if (cs==READY) begin
    end

end


//////////////////////////////////



endmodule
